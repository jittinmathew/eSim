* C:\Users\Jittin\eSim-Workspace\RC\RC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 08/26/21 10:15:20

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  OUT IN 1k		
C1  OUT GND 1u		
v1  IN GND sine		
U2  OUT plot_v1		
U1  IN plot_v1		

.end
